module MEM_WB_Reg (
    input wire clk,
    input wire rst,

    input wire [1:0] mem_to_reg_i,
    input wire regWrite_i,
    input wire [31:0] pc_4_i,
    input wire [4:0] writeReg_i,
    input wire [31:0] ALU_result_i,
    input wire [31:0] readDataResult_i,

    output reg [1:0] mem_to_reg_o,
    output reg regWrite_o,
    output reg [31:0] pc_4_o,
    output reg [4:0] writeReg_o,
    output reg [31:0] ALU_result_o,
    output reg [31:0] readDataResult_o
);

    always @(posedge clk or negedge rst) begin
        if (~rst) begin
            mem_to_reg_o <= mem_to_reg_o;
            regWrite_o <= regWrite_o;
            pc_4_o <= pc_4_o;
            writeReg_o <= writeReg_o;
            ALU_result_o <= ALU_result_o;
            readDataResult_o <= readDataResult_o;
        end 
        else begin
            mem_to_reg_o <= mem_to_reg_i;
            regWrite_o <= regWrite_i;
            pc_4_o <= pc_4_i;
            writeReg_o <= writeReg_i;
            ALU_result_o <= ALU_result_i;
            readDataResult_o <= readDataResult_i;
        end
    end

endmodule
